module Divisor (
    input [31:0] Dvsr_in,
    output [31:0] Dvsr_out
);
    assign Dvsr_out = Dvsr_in;
endmodule