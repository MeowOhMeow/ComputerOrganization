module Multiplicand (
    input [31:0] Mult_in,
    output [31:0] Mult_out
);
    assign Mult_out = Mult_in;

endmodule